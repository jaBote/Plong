library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity bar_rom is
    port(
        clk: in std_logic;
        addr: in std_logic_vector(5 downto 0);
        data: out std_logic_vector(0 to 127)
    );
end bar_rom;

architecture content of bar_rom is
    type rom_type is array(0 to 19) of std_logic_vector(127 downto 0);
    constant BAR: rom_type :=
    (
		"11111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111101111111111110",
		"11000000000000010000010000000100000000001000010100010000001000001010000000000000000000000010100010101010100000000010000010001010",
		"10101111111101101111010111111011111111110101010111101011110100110010101111111110111011101001011011011001011111101101111010110110",
		"11110000000000000000000000001110000000000000000001010100001000001000000000000000000100000000100001111110100000000000000000001010",
		"10011110100010110000000000100101111000000000000000010000110101010100000001000000100010010110011111101011110100010110000000000110",
		"11000111101100000000000000011101000000000000001000000101000010101010000110100000000000001001101110000000111101100000000000001110",
		"00100001110001010000101100101100000000000010010010110100110000000000000000000000000011100111100000000000001110001010000101100010",
		"10000000011010000000000011011000010001000000000001000111001101001001101010000000000000111110000000000000000011010000000000011110",
		"10110000000100001000100000110010000000000000000000000001110010100110000100011000000001111000000000000001000000100001000100000110",
		"10000000011010110010001011100000000000000011001000001101011100010000100000000000010111100000000000000010000011010110010001011110",
		"10100011000101001000110100110000000000000000010000000000000101011110000000000000001010000001000000010000011000101001000110101110",
		"10000000100011101101001011000000100000001000000101011100010100100000000000000000010110000000000000100100000100011101101001011010",
		"10110000000100111010111100000000010001000000000000000000000000000110001000000001011110000000000000001001000000100111010111100110",
		"10000000110000000101110000000011000000110000000000110010000000000000000110000110101100000000011000000010000110000000101110001010",
		"10100000001100101011000011001100000000000000000010000000001000011100010000001001110000000100000001000000000001100101011000010110",
		"11001000010000010100000000010000001011000000001001101100100000100100001010010111000000011000000100000001000010000010100000001010",
		"00100000100000000000000000000010000000000000000000000000101000011111100001101100000001000000000001000000000100000000000000000110",
		"10110111011111001010101010101001111101110010101010110010100111000000010101011001011001010101010100010110111011111001010101011110",
		"10001000100000101010101010101010000010001010101011001010101000111101111111110101000101010101010101010001000100000101010101010110",
		"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"
    );
    signal addr_reg: std_logic_vector(5 downto 0);
begin
    process(clk)
    begin
        if clk'event and clk = '1' then
            addr_reg <= addr;
        end if;
    end process;            
    data <= BAR(conv_integer(addr_reg));
end content;

