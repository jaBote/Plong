library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity brick_rom is
    port(
        addr: in std_logic_vector(4 downto 0);
        data: out std_logic_vector(0 to 39)
    );
end brick_rom;

architecture content of brick_rom is
    type rom_type is array(0 to 19) of std_logic_vector(39 downto 0);
    constant BRICK: rom_type :=
    (
        "1111111111111111111111111111111111111111",
        "1011000000000000000000000000000000001101",
        "1000110000000000000000000000000000110001",
        "1000001100000000000000000000000011000001",
        "1000000011000000000000000000001100000001",
        "1000000000110000000000000000110000000001",
        "1000000000001100000000000011000000000001",
        "1000000000000011000000001100000000000001",
        "1000000000000000110000110000000000000001",
        "1000000000000000001111000000000000000001",
        "1000000000000000001111000000000000000001",
        "1000000000000000110000110000000000000001",
        "1000000000000011000000001100000000000001",
        "1000000000001100000000000011000000000001",
        "1000000000110000000000000000110000000001",
        "1000000011000000000000000000001100000001",
        "1000001100000000000000000000000011000001",
        "1000110000000000000000000000000000110001",
        "1011000000000000000000000000000000001101",
        "1111111111111111111111111111111111111111"
    );
begin
    data <= BRICK(conv_integer(addr));
end content;
